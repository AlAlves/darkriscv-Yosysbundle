module rvfi_wrapper (
	input clock,
	input reset,
	`RVFI_OUTPUTS
);


	darkriscv uut (

	)





endmodule
